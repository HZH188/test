module leg (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input;
  output  wire [7:0] Output;

  TC_Register # (.UUID(64'd948720666095222483 ^ UUID), .BIT_WIDTH(64'd8)) Register8_0 (.clk(clk), .rst(rst), .load(wire_8), .save(wire_47), .in(wire_44), .out(wire_34));
  TC_Register # (.UUID(64'd3288173254724515669 ^ UUID), .BIT_WIDTH(64'd8)) Register8_1 (.clk(clk), .rst(rst), .load(wire_92), .save(wire_11), .in(wire_79), .out(wire_12));
  TC_Register # (.UUID(64'd2138514348962238939 ^ UUID), .BIT_WIDTH(64'd8)) Register8_2 (.clk(clk), .rst(rst), .load(wire_57), .save(wire_81), .in(wire_29), .out(wire_40));
  TC_Register # (.UUID(64'd2719339641550232870 ^ UUID), .BIT_WIDTH(64'd8)) Register8_3 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_74), .in(wire_77), .out(wire_70));
  TC_Register # (.UUID(64'd1118205527678439814 ^ UUID), .BIT_WIDTH(64'd8)) Register8_4 (.clk(clk), .rst(rst), .load(wire_93), .save(wire_48), .in(wire_96), .out(wire_51));
  TC_Switch # (.UUID(64'd2465942727236428333 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_47), .in(wire_17), .out(wire_44));
  TC_Switch # (.UUID(64'd1566235650929549540 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_11), .in(wire_17), .out(wire_79));
  TC_Switch # (.UUID(64'd3449418223612905723 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_81), .in(wire_17), .out(wire_29));
  TC_Switch # (.UUID(64'd99626139207926688 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_74), .in(wire_17), .out(wire_77));
  TC_Switch # (.UUID(64'd3914604852771176598 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_48), .in(wire_17), .out(wire_96));
  TC_Switch # (.UUID(64'd712410099928060352 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_30), .in(wire_17), .out(wire_97));
  TC_Switch # (.UUID(64'd795442694490214132 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_42), .in(wire_34), .out(wire_3_0));
  TC_Switch # (.UUID(64'd1423286731315913415 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_41), .in(wire_12), .out(wire_3_1));
  TC_Switch # (.UUID(64'd314329153825463881 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_23), .in(wire_40), .out(wire_3_2));
  TC_Switch # (.UUID(64'd4305714527704135472 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_88), .in(wire_70), .out(wire_3_3));
  TC_Switch # (.UUID(64'd355662053832162974 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_28), .in(wire_51), .out(wire_3_4));
  TC_Switch # (.UUID(64'd2686953195933991358 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_78), .in(wire_83), .out(wire_3_6));
  TC_Constant # (.UUID(64'd4248611437735476737 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out(wire_8));
  TC_Constant # (.UUID(64'd62872831037185520 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_18 (.out(wire_92));
  TC_Constant # (.UUID(64'd868267106323219813 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_19 (.out(wire_57));
  TC_Constant # (.UUID(64'd4567596755233995393 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_20 (.out(wire_24));
  TC_Constant # (.UUID(64'd1983339691876125001 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_21 (.out(wire_93));
  TC_Constant # (.UUID(64'd3681301743804406468 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_22 (.out(wire_98));
  TC_Register # (.UUID(64'd1103605438749734585 ^ UUID), .BIT_WIDTH(64'd8)) Register8_23 (.clk(clk), .rst(rst), .load(wire_98), .save(wire_30), .in(wire_97), .out(wire_83));
  TC_Switch # (.UUID(64'd2742420798102234718 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_46), .in(wire_6), .out(wire_25_8));
  TC_Switch # (.UUID(64'd3615289143049369418 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_55), .in(wire_17), .out(wire_49));
  TC_Splitter8 # (.UUID(64'd1973025975119237032 ^ UUID)) Splitter8_26 (.in({{7{1'b0}}, wire_2 }), .out0(wire_33), .out1(wire_76), .out2(wire_10), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd241159497683819979 ^ UUID)) Decoder3_27 (.dis(wire_94), .sel0(wire_33), .sel1(wire_76), .sel2(wire_10), .out0(wire_1), .out1(wire_52), .out2(wire_80), .out3(wire_108), .out4(wire_71), .out5(wire_68), .out6(wire_62), .out7(wire_46));
  TC_Splitter8 # (.UUID(64'd112032136428255408 ^ UUID)) Splitter8_28 (.in({{7{1'b0}}, wire_36 }), .out0(wire_117), .out1(wire_67), .out2(wire_61), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2903030717399396891 ^ UUID)) Decoder3_29 (.dis(wire_114), .sel0(wire_117), .sel1(wire_67), .sel2(wire_61), .out0(wire_42), .out1(wire_41), .out2(wire_23), .out3(wire_88), .out4(wire_28), .out5(wire_78), .out6(wire_26), .out7(wire_27));
  TC_Splitter8 # (.UUID(64'd3434298155437954163 ^ UUID)) Splitter8_30 (.in({{7{1'b0}}, wire_31 }), .out0(wire_65), .out1(wire_118), .out2(wire_116), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd2584112576133784572 ^ UUID)) Decoder3_31 (.dis(wire_60), .sel0(wire_65), .sel1(wire_118), .sel2(wire_116), .out0(wire_47), .out1(wire_11), .out2(wire_81), .out3(wire_74), .out4(wire_48), .out5(wire_30), .out6(wire_4), .out7(wire_55));
  TC_Switch # (.UUID(64'd2968724590403814568 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_32 (.en(wire_27), .in(wire_6), .out(wire_3_8));
  TC_Switch # (.UUID(64'd852776023643561415 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_1), .in(wire_34), .out(wire_25_0));
  TC_Switch # (.UUID(64'd2811511616213636218 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_34 (.en(wire_52), .in(wire_12), .out(wire_25_1));
  TC_Switch # (.UUID(64'd4336349970457983445 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_35 (.en(wire_80), .in(wire_40), .out(wire_25_2));
  TC_Switch # (.UUID(64'd2387349439961323536 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_36 (.en(wire_108), .in(wire_70), .out(wire_25_4));
  TC_Switch # (.UUID(64'd2424276507761906001 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_37 (.en(wire_71), .in(wire_51), .out(wire_25_6));
  TC_Switch # (.UUID(64'd439621575481776013 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_38 (.en(wire_68), .in(wire_83), .out(wire_25_7));
  TC_Constant # (.UUID(64'd2657984117251512804 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_39 (.out(wire_113));
  TC_Splitter8 # (.UUID(64'd4300721551118231460 ^ UUID)) Splitter8_40 (.in(wire_0), .out0(wire_7), .out1(wire_22), .out2(wire_99), .out3(wire_90), .out4(wire_111), .out5(wire_63), .out6(wire_13), .out7(wire_66));
  TC_Maker8 # (.UUID(64'd143746129312731296 ^ UUID)) Maker8_41 (.in0(wire_7), .in1(wire_22), .in2(wire_99), .in3(wire_90), .in4(wire_111), .in5(wire_63), .in6(wire_13), .in7(wire_66), .out(wire_86));
  TC_Switch # (.UUID(64'd1857701737722394134 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_42 (.en(wire_66), .in({{7{1'b0}}, wire_2 }), .out(wire_25_3));
  TC_Not # (.UUID(64'd2439651504842858841 ^ UUID), .BIT_WIDTH(64'd1)) Not_43 (.in(1'd0), .out(wire_43));
  TC_Switch # (.UUID(64'd2909453999051889468 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_43), .in(wire_59), .out(wire_17));
  TC_Equal # (.UUID(64'd3685796226974449157 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_45 (.in0(wire_109), .in1(wire_39), .out(wire_56));
  TC_Switch # (.UUID(64'd1004915224443871815 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_46 (.en(wire_20[0:0]), .in(wire_25), .out(wire_109));
  TC_Switch # (.UUID(64'd1966495235752351639 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_20[0:0]), .in(wire_3), .out(wire_39));
  TC_Switch # (.UUID(64'd1597509329047381879 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_38[0:0]), .in(wire_25), .out(wire_89));
  TC_Equal # (.UUID(64'd2833496657859985473 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_49 (.in0(wire_89), .in1(wire_91), .out(wire_73));
  TC_Switch # (.UUID(64'd852619902536349452 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_38[0:0]), .in(wire_3), .out(wire_91));
  TC_Switch # (.UUID(64'd2937067025135784017 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_51 (.en(wire_20[0:0]), .in(wire_56), .out(wire_15_5));
  TC_Switch # (.UUID(64'd2936443805849482296 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_52 (.en(wire_38[0:0]), .in(wire_50), .out(wire_15_4));
  TC_Not # (.UUID(64'd2348731379215183627 ^ UUID), .BIT_WIDTH(64'd1)) Not_53 (.in(wire_73), .out(wire_50));
  TC_Switch # (.UUID(64'd3448084879071483539 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_19[0:0]), .in(wire_25), .out(wire_69));
  TC_Switch # (.UUID(64'd1979956127529990309 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_55 (.en(wire_19[0:0]), .in(wire_3), .out(wire_85));
  TC_Switch # (.UUID(64'd4541042300876392443 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_56 (.en(wire_19[0:0]), .in(wire_101), .out(wire_15_3));
  TC_LessU # (.UUID(64'd493087175006901653 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_57 (.in0(wire_69), .in1(wire_85), .out(wire_101));
  TC_LessU # (.UUID(64'd1859070900694287058 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_58 (.in0(wire_105), .in1(wire_87), .out(wire_9));
  TC_Switch # (.UUID(64'd1490513829384869263 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_59 (.en(wire_16[0:0]), .in(wire_25), .out(wire_105));
  TC_Switch # (.UUID(64'd873754934868526673 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_60 (.en(wire_16[0:0]), .in(wire_3), .out(wire_87));
  TC_Switch # (.UUID(64'd676521216694563762 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_61 (.en(wire_16[0:0]), .in(wire_82), .out(wire_15_0));
  TC_Not # (.UUID(64'd760413059066947120 ^ UUID), .BIT_WIDTH(64'd1)) Not_62 (.in(wire_9), .out(wire_82));
  TC_Switch # (.UUID(64'd1328255739527756627 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_63 (.en(wire_43), .in({{7{1'b0}}, wire_37 }), .out(wire_0));
  TC_Switch # (.UUID(64'd2898445796686407799 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_64 (.en(wire_54[0:0]), .in(wire_25), .out(wire_115));
  TC_Switch # (.UUID(64'd1081244702047706055 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_65 (.en(wire_54[0:0]), .in(wire_3), .out(wire_84));
  TC_Switch # (.UUID(64'd1399805028219565247 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_66 (.en(wire_54[0:0]), .in(wire_18[0:0]), .out(wire_15_1));
  TC_Switch # (.UUID(64'd131407806234628885 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_67 (.en(wire_21[0:0]), .in(wire_25), .out(wire_112));
  TC_Switch # (.UUID(64'd449638382667490273 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_68 (.en(wire_21[0:0]), .in(wire_3), .out(wire_107));
  TC_Switch # (.UUID(64'd1328437419064840760 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_69 (.en(wire_21[0:0]), .in(wire_95), .out(wire_15_2));
  TC_Not # (.UUID(64'd2207909349942323425 ^ UUID), .BIT_WIDTH(64'd1)) Not_70 (.in(wire_100[0:0]), .out(wire_95));
  TC_Switch # (.UUID(64'd1733094870635544701 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_71 (.en(wire_13), .in({{7{1'b0}}, wire_36 }), .out(wire_3_7));
  TC_Switch # (.UUID(64'd4196173604070654814 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_72 (.en(wire_4), .in(wire_17), .out(wire_53_2));
  TC_Counter # (.UUID(64'd3477379483004833537 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_73 (.clk(clk), .rst(rst), .save(wire_106), .in(wire_53), .out(wire_14));
  TC_Switch # (.UUID(64'd556936333953868570 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_74 (.en(wire_102), .in({{7{1'b0}}, wire_31 }), .out(wire_53_0));
  TC_Switch # (.UUID(64'd2561998164344676762 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_62), .in(wire_14), .out(wire_25_5));
  TC_Switch # (.UUID(64'd1014432617426286536 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_76 (.en(wire_26), .in(wire_14), .out(wire_3_5));
  TC_Constant # (.UUID(64'd1550467710238502600 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_77 (.out(wire_110));
  TC_Equal # (.UUID(64'd4527919892871818404 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_78 (.in0({{7{1'b0}}, wire_37 }), .in1(wire_110), .out(wire_45));
  TC_Add # (.UUID(64'd2933028734573733631 ^ UUID), .BIT_WIDTH(64'd8)) Add8_79 (.in0(wire_14), .in1(wire_103), .ci(1'd0), .out(wire_104), .co());
  TC_Constant # (.UUID(64'd3972693244687706560 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_80 (.out(wire_103));
  TC_Or # (.UUID(64'd1782278601304283403 ^ UUID), .BIT_WIDTH(64'd1)) Or_81 (.in0(wire_45), .in1(wire_15), .out(wire_102));
  TC_Equal # (.UUID(64'd1169725261175755572 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_82 (.in0({{7{1'b0}}, wire_37 }), .in1(wire_72), .out(wire_5));
  TC_Constant # (.UUID(64'd115174148557746969 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h10)) Constant8_83 (.out(wire_72));
  TC_Switch # (.UUID(64'd1256829898421007229 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_84 (.en(wire_5), .in(wire_64), .out(wire_53_1));
  TC_Or3 # (.UUID(64'd1903221479974050264 ^ UUID), .BIT_WIDTH(64'd1)) Or3_85 (.in0(wire_15), .in1(wire_58), .in2(wire_4), .out(wire_106));
  TC_Or # (.UUID(64'd1653749908697703264 ^ UUID), .BIT_WIDTH(64'd1)) Or_86 (.in0(wire_5), .in1(wire_45), .out(wire_58));
  TC_Or # (.UUID(64'd770855609776920846 ^ UUID), .BIT_WIDTH(64'd1)) Or_87 (.in0(wire_35[0:0]), .in1(wire_58), .out(wire_60));
  TC_Or # (.UUID(64'd760423012748264367 ^ UUID), .BIT_WIDTH(64'd1)) Or_88 (.in0(wire_13), .in1(wire_32[0:0]), .out(wire_114));
  TC_Or # (.UUID(64'd1371424513914838714 ^ UUID), .BIT_WIDTH(64'd1)) Or_89 (.in0(wire_66), .in1(wire_75[0:0]), .out(wire_94));
  greaterz_than # (.UUID(64'd2345821357778772423 ^ UUID)) greaterz_than_90 (.clk(clk), .rst(rst), .Input_1(wire_112), .Input_2(wire_107), .Output(wire_100));
  calcuate2 # (.UUID(64'd779880426580832613 ^ UUID)) calcuate2_91 (.clk(clk), .rst(rst), .\�_____ (wire_86), .\�______1 (wire_25), .\�______2 (wire_3), .Output(wire_59));
  greaterz_than # (.UUID(64'd4496997152499601284 ^ UUID)) greaterz_than_92 (.clk(clk), .rst(rst), .Input_1(wire_115), .Input_2(wire_84), .Output(wire_18));
  ZXE6ZXA0ZX88 # (.UUID(64'd1906505505157829066 ^ UUID)) ZXE6ZXA0ZX88_93 (.clk(clk), .rst(rst), .POP(wire_5), .PUSH(wire_45), .VALUE(wire_104), .OUTPUT(wire_64));
  choosez_3 # (.UUID(64'd3590042652547995650 ^ UUID)) choosez_3_94 (.clk(clk), .rst(rst), .Input({{7{1'b0}}, wire_37 }), .Output_1(wire_20), .Output_2(wire_38), .Output_3(wire_19), .Output_4(wire_21), .Output_5(wire_54), .Output_6(wire_16), .Output_7(wire_35));
  lock # (.UUID(64'd948675432539824519 ^ UUID)) lock_95 (.clk(clk), .rst(rst), .Input_1({{7{1'b0}}, wire_36 }), .Input_2({{7{1'b0}}, wire_2 }), .Output_1(wire_32), .Output_2(wire_75));

  wire [7:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  assign wire_2 = 0;
  wire [7:0] wire_3;
  wire [7:0] wire_3_0;
  wire [7:0] wire_3_1;
  wire [7:0] wire_3_2;
  wire [7:0] wire_3_3;
  wire [7:0] wire_3_4;
  wire [7:0] wire_3_5;
  wire [7:0] wire_3_6;
  wire [7:0] wire_3_7;
  wire [7:0] wire_3_8;
  assign wire_3 = wire_3_0|wire_3_1|wire_3_2|wire_3_3|wire_3_4|wire_3_5|wire_3_6|wire_3_7|wire_3_8;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  assign wire_6 = Input;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_15_0;
  wire [0:0] wire_15_1;
  wire [0:0] wire_15_2;
  wire [0:0] wire_15_3;
  wire [0:0] wire_15_4;
  wire [0:0] wire_15_5;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2|wire_15_3|wire_15_4|wire_15_5;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_25_0;
  wire [7:0] wire_25_1;
  wire [7:0] wire_25_2;
  wire [7:0] wire_25_3;
  wire [7:0] wire_25_4;
  wire [7:0] wire_25_5;
  wire [7:0] wire_25_6;
  wire [7:0] wire_25_7;
  wire [7:0] wire_25_8;
  assign wire_25 = wire_25_0|wire_25_1|wire_25_2|wire_25_3|wire_25_4|wire_25_5|wire_25_6|wire_25_7|wire_25_8;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [7:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  assign wire_31 = 0;
  wire [7:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  assign wire_36 = 0;
  wire [0:0] wire_37;
  assign wire_37 = 0;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [7:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [7:0] wire_49;
  assign Output = wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [7:0] wire_53;
  wire [7:0] wire_53_0;
  wire [7:0] wire_53_1;
  wire [7:0] wire_53_2;
  assign wire_53 = wire_53_0|wire_53_1|wire_53_2;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [7:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [7:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [7:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [7:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [7:0] wire_77;
  wire [0:0] wire_78;
  wire [7:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [7:0] wire_83;
  wire [7:0] wire_84;
  wire [7:0] wire_85;
  wire [7:0] wire_86;
  wire [7:0] wire_87;
  wire [0:0] wire_88;
  wire [7:0] wire_89;
  wire [0:0] wire_90;
  wire [7:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [7:0] wire_96;
  wire [7:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [7:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [7:0] wire_103;
  wire [7:0] wire_104;
  wire [7:0] wire_105;
  wire [0:0] wire_106;
  wire [7:0] wire_107;
  wire [0:0] wire_108;
  wire [7:0] wire_109;
  wire [7:0] wire_110;
  wire [0:0] wire_111;
  wire [7:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [7:0] wire_115;
  wire [0:0] wire_116;
  wire [0:0] wire_117;
  wire [0:0] wire_118;

endmodule
